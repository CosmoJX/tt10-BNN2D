`include "Conv2d.sv"
`include "MaxPool2d.sv"

module dut (
    // input logic [CONV1_IMG_IN_SIZE*CONV1_IMG_IN_SIZE-1:0] img_in [0:CONV1_IC-1]
);
    parameter int CONV1_IC = 1;
    parameter int CONV1_OC = 10;
    parameter int CONV2_OC = 8;
    parameter int FC_IC= POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE*CONV2_OC;
    parameter int FC_OC = 10;                   // num classes
    parameter int CONV1_IMG_IN_SIZE = 30;
    parameter int CONV1_IMG_OUT_SIZE = CONV1_IMG_IN_SIZE-2;
    parameter int POOL1_IMG_OUT_SIZE = CONV1_IMG_OUT_SIZE/2;
    parameter int CONV2_IMG_OUT_SIZE = POOL1_IMG_OUT_SIZE-2;
    parameter int POOL2_IMG_OUT_SIZE = CONV2_IMG_OUT_SIZE/2;
    parameter int OUTPUT_BIT = $clog2(FC_OC+1); // num of bits to enumerate each class

    logic [CONV1_IMG_IN_SIZE*CONV1_IMG_IN_SIZE-1:0] conv1_img_in [0:CONV1_IC-1] = {900'h1e000000ff000003fe00000c38000030700000c1c00003f7000007fc000007f0000001c000000700000038000001e000000f000000f8000003c000000c000000000000000000000000000000000000000000000000000000000};
    // assign conv1_img_in = img_in;
    logic [CONV1_IC*9-1:0] conv1_weights [0:CONV1_OC-1] = {9'hde, 9'h183, 9'h98, 9'h3e, 9'h1d6, 9'h6e, 9'h17c, 9'hf9, 9'hc9, 9'h18a};
    logic [CONV1_OC*9-1:0] conv2_weights [0:CONV2_OC-1] = {90'h1eecfbdb3c7b7800819e, 90'h224e92fb00d30024868, 90'h5a00381c70144e800003d, 90'h882d020940a259200179, 90'hb8e07048ff6638000182, 90'h2ffcda1933be868401a8, 90'he1b86120106c28800b0, 90'hf4e1b0881d2e444001b6};
    logic signed [15:0] fc_weights [0:FC_IC*FC_OC-1] = {16'hfffb, 16'h10, 16'h6, 16'h47, 16'h1e, 16'h0, 16'hffef, 16'hffe3, 16'hffce, 16'hffcb, 16'h2, 16'hfffc, 
                                                     16'hffe2, 16'hff8f, 16'hff9d, 16'hffbb, 16'hff97, 16'h0, 16'hffea, 16'hffc2, 16'hff99, 16'hff6c, 16'hff4a, 
                                                     16'hffed, 16'hffe3, 16'h25, 16'hffa0, 16'hff79, 16'hffa9, 16'hffee, 16'hffe8, 16'h4a, 16'h30, 16'h3b, 16'h26, 
                                                     16'h1b, 16'h3, 16'hffdd, 16'h1d, 16'h12, 16'hffcd, 16'hfff8, 16'ha, 16'h7, 16'h14, 16'hb9, 16'h88, 16'h4, 16'h68, 
                                                     16'h49, 16'h94, 16'he8, 16'h11d, 16'h6, 16'hb8, 16'ha6, 16'hab, 16'hee, 16'hf9, 16'h2a, 16'h6e, 16'h67, 16'h42, 
                                                     16'h4b, 16'h65, 16'hfff2, 16'h37, 16'h13, 16'hffc0, 16'hffa4, 16'hff80, 16'hffe8, 16'h39, 16'h21, 16'hffe6, 
                                                     16'hffe6, 16'hffea, 16'h1b, 16'h20, 16'hffb0, 16'hff6a, 16'hffb2, 16'hffe6, 16'hffe7, 16'h1b, 16'hff5b, 16'hff2f, 
                                                     16'hff42, 16'hff9c, 16'hffcd, 16'hffcb, 16'hff6e, 16'hff70, 16'hff99, 16'hffe7, 16'hffee, 16'hffee, 16'hfffb, 
                                                     16'hfff4, 16'hfff6, 16'h9, 16'hfffc, 16'h0, 16'hc, 16'h12, 16'h1c, 16'h16, 16'h5, 16'h12, 16'h1c, 16'hffc7, 16'hffe2, 
                                                     16'hffc2, 16'hffb1, 16'hfffe, 16'h1d, 16'h7a, 16'hffda, 16'hff83, 16'hffac, 16'hffd9, 16'h60, 16'hae, 16'hffef, 
                                                     16'hfffa, 16'h19, 16'hffda, 16'h84, 16'h8b, 16'h6b, 16'h68, 16'h55, 16'hffd3, 16'h10, 16'h4, 16'h1c, 16'h4b, 16'h44, 
                                                     16'h2, 16'hffdf, 16'hffc7, 16'hffd0, 16'h34, 16'h41, 16'hffed, 16'hffc5, 16'h8, 16'h21, 16'hffdf, 16'hffdc, 16'hffd6, 
                                                     16'h9, 16'h1a, 16'h29, 16'hffca, 16'hffd8, 16'h1, 16'hffea, 16'hffa3, 16'hff84, 16'hffa1, 16'hffd5, 16'hffdb, 
                                                     16'hffa0, 16'hff78, 16'hff71, 16'hffb3, 16'hffc4, 16'hfff2, 16'hffd8, 16'hffdf, 16'hffd1, 16'hfffa, 16'hffe5, 
                                                     16'hfff2, 16'hffe5, 16'h13, 16'h16, 16'he, 16'hfff5, 16'h11, 16'h14, 16'h31, 16'h53, 16'h1d, 16'h6, 16'h22, 
                                                     16'hffeb, 16'hd, 16'h4a, 16'h28, 16'h27, 16'h1b, 16'h2f, 16'h17, 16'h10, 16'h25, 16'h23, 16'hfff3, 16'h18, 16'h18, 16'h0, 
                                                     16'h1a, 16'h1a, 16'h3, 16'h17, 16'h52, 16'h1d, 16'hfff8, 16'hffe3, 16'h3, 16'h22, 16'h50, 16'h44, 16'h2d, 16'hfffe, 16'h2b, 
                                                     16'h31, 16'hffd0, 16'hffb1, 16'hffe5, 16'h14, 16'h3a, 16'hfff9, 16'hfff1, 16'hffa8, 16'hffc9, 16'hffd8, 16'h33, 16'hffcc, 
                                                     16'hff90, 16'hff8e, 16'hffa8, 16'hff96, 16'hfffb, 16'hff93, 16'hff97, 16'h4, 16'hffec, 16'hffc1, 16'hffe2, 16'hffc3, 16'hffe0, 
                                                     16'hfff7, 16'hfffb, 16'hffdf, 16'hffef, 16'hffe5, 16'hffe9, 16'hffeb, 16'hfffc, 16'h21, 16'hffdf, 16'hffd5, 16'hfffa, 16'h2e, 
                                                     16'hffe3, 16'h6, 16'hfff0, 16'h3, 16'hfffb, 16'h46, 16'hfffb, 16'h17, 16'h24, 16'h47, 16'h58, 16'h32, 16'h38, 16'h53, 16'h7, 
                                                     16'h6c, 16'h5a, 16'h2c, 16'h36, 16'h34, 16'hc, 16'h3a, 16'h46, 16'h2b, 16'h19, 16'hc, 16'he, 16'h20, 16'h21, 16'h15, 16'h11, 
                                                     16'hfff9, 16'h39, 16'h50, 16'hffd6, 16'hff6c, 16'hffc3, 16'h3d, 16'h6e, 16'h26, 16'hff48, 16'hff82, 16'hffc8, 16'hf, 16'h4e, 
                                                     16'hffe1, 16'hff74, 16'hffc4, 16'hffdf, 16'hffe0, 16'h4d, 16'hff9c, 16'hff68, 16'hffbb, 16'hffc0, 16'hd, 16'h5b, 16'hffd7, 
                                                     16'hff7a, 16'hff7b, 16'hffbe, 16'h3, 16'h2f, 16'hc, 16'hffbc, 16'hffb6, 16'hffea, 16'h6, 16'h3a, 16'hffd0, 16'h3f, 16'h81, 
                                                     16'h59, 16'h3b, 16'h2, 16'hffe5, 16'h69, 16'h83, 16'h30, 16'h64, 16'hffc9, 16'hfff2, 16'h51, 16'h56, 16'h14, 16'h58, 16'hffc0, 
                                                     16'h14, 16'h39, 16'h6f, 16'hc, 16'h54, 16'h19, 16'h5b, 16'h73, 16'h9a, 16'h2f, 16'h42, 16'hd, 16'h21, 16'h72, 16'h88, 16'h5c, 
                                                     16'h70, 16'h45, 16'h55, 16'h63, 16'h6d, 16'h71, 16'h1e, 16'h3c, 16'h16, 16'hffe5, 16'h29, 16'h5f, 16'h46, 16'h2b, 16'hffe7, 
                                                     16'hfffd, 16'h1d, 16'h1e, 16'h61, 16'hffde, 16'hffb8, 16'hffc7, 16'hfff8, 16'hd, 16'h1b, 16'h7, 16'hffc8, 16'hffa7, 16'hffbe, 
                                                     16'hb, 16'h7, 16'h1e, 16'hffdf, 16'hffb9, 16'hffc8, 16'hffe9, 16'h3, 16'h61, 16'h69, 16'h7a, 16'h30, 16'hffcf, 16'hffd2, 16'h53, 
                                                     16'h4c, 16'hc2, 16'h33, 16'hffd6, 16'hffb8, 16'h5c, 16'h5b, 16'hc9, 16'h16, 16'hffe5, 16'hffcb, 16'h4c, 16'h3f, 16'h5e, 16'hfff6, 
                                                     16'hffed, 16'hffa2, 16'h34, 16'h79, 16'h83, 16'h54, 16'h21, 16'hffdd, 16'h64, 16'h86, 16'h60, 16'h40, 16'h1c, 16'hffd8, 16'h5a, 
                                                     16'hfffe, 16'hffa7, 16'hffd3, 16'hffed, 16'h1, 16'h41, 16'hffe6, 16'hff96, 16'hffb3, 16'hffcb, 16'hffea, 16'h30, 16'hffd7, 16'hffa5, 
                                                     16'hffb5, 16'hffbd, 16'hffe6, 16'h2e, 16'hffea, 16'hffa3, 16'hff9d, 16'hffb7, 16'hfff9, 16'h47, 16'hfff9, 16'hffdf, 16'hffba, 16'hffeb, 
                                                     16'hc, 16'h60, 16'h30, 16'h1a, 16'hfff8, 16'h18, 16'h33, 16'hfffd, 16'hff77, 16'hff8e, 16'hff79, 16'hff7d, 16'hffbc, 16'hfff0, 16'hffa2, 
                                                     16'hff8f, 16'hff8a, 16'hff95, 16'hffcd, 16'hffbe, 16'hff6e, 16'hff65, 16'hff64, 16'hff72, 16'hffce, 16'hffc6, 16'hff89, 16'hff4e, 16'hff6c, 
                                                     16'hff5e, 16'hffd2, 16'hffec, 16'hffc5, 16'hffa0, 16'hffb9, 16'hffa4, 16'hffe0, 16'h21, 16'hffdd, 16'hffc8, 16'hffcc, 16'hffe9, 16'hffd0, 
                                                     16'hffbd, 16'hffd3, 16'h62, 16'h7f, 16'h34, 16'hffe8, 16'hffc2, 16'hfff6, 16'h4c, 16'h42, 16'h37, 16'h25, 16'hffd2, 16'h26, 16'h4a, 16'h25, 
                                                     16'h2e, 16'h14, 16'hffec, 16'h3a, 16'h4, 16'h8, 16'hfffc, 16'h17, 16'hffe0, 16'h26, 16'h33, 16'h23, 16'h1a, 16'hfffa, 16'hffda, 16'h4, 
                                                     16'h30, 16'h1f, 16'h16, 16'hfff0, 16'h2a, 16'hffba, 16'hff9b, 16'hffba, 16'hffd3, 16'hffa6, 16'h68, 16'hff8f, 16'hff76, 16'hffb8, 16'hffd6, 
                                                     16'hff83, 16'h9, 16'hff8b, 16'hffba, 16'hffd6, 16'hffb7, 16'hff92, 16'h27, 16'hffbe, 16'hffc9, 16'hffc1, 16'hffd3, 16'hffbd, 16'h35, 16'hfff0, 
                                                     16'h2, 16'hffed, 16'hffe7, 16'hffe2, 16'h52, 16'h11, 16'h7, 16'h3, 16'hfff2, 16'hffdd, 16'hffb9, 16'hffb0, 16'hff9d, 16'hffb2, 16'hffce, 
                                                     16'hffdc, 16'hffd9, 16'hffc4, 16'hff6e, 16'hff5e, 16'hffb3, 16'hffca, 16'hffc3, 16'hff85, 16'hff6d, 16'hff5b, 16'hff84, 16'hffbb, 16'hffdf, 
                                                     16'hffbd, 16'hffa4, 16'hffbb, 16'hffdb, 16'h3, 16'hffe9, 16'hffd2, 16'h6, 16'h3b, 16'h55, 16'h2c, 16'hffec, 16'hffe5, 16'h5c, 16'h9f, 16'h43, 
                                                     16'h17, 16'hffd9, 16'hffd1, 16'hffef, 16'hffb4, 16'hffd0, 16'hffcd, 16'hffb9, 16'hffdb, 16'hffbf, 16'h26, 16'h2e, 16'hffdf, 16'hff6d, 16'hff7e, 
                                                     16'hffb0, 16'h59, 16'h7f, 16'hffeb, 16'hffa4, 16'hff77, 16'hff87, 16'h1, 16'h12, 16'hffe3, 16'hffe0, 16'hffc1, 16'hff8b, 16'hff49, 16'hff3e, 
                                                     16'hffd7, 16'hfff2, 16'hffba, 16'hffaa, 16'hff47, 16'hffac, 16'hffd4, 16'hffa8, 16'hffad, 16'hffe2, 16'hffc6, 16'hffc3, 16'hffd7, 16'hffac, 
                                                     16'hbb, 16'h104, 16'h60, 16'h7, 16'hffb7, 16'hffb5, 16'h54, 16'hae, 16'h73, 16'h2e, 16'hffdb, 16'h58, 16'hc6, 16'hc6, 16'hc2, 16'hdd, 16'h99, 
                                                     16'h5f, 16'h7f, 16'h8f, 16'hba, 16'hbb, 16'haa, 16'h21, 16'h33, 16'h75, 16'hb5, 16'h85, 16'h54, 16'hffec, 16'hfff1, 16'hffd8, 16'hffa4, 16'hff45, 16'hff85, 16'hffd3, 16'hffd5, 16'h2, 16'hffdf, 16'hffa5, 16'hffba, 16'hffdb, 16'hff9a, 16'h13, 16'hfff5, 16'h6, 16'h1c, 16'hffb5, 16'h75, 16'h5f, 16'hfff6, 16'hffff, 16'hb, 16'hffd5, 16'h6b, 16'h48, 16'hffc9, 16'hffbd, 16'hffcd, 16'hffdc, 16'h53, 16'h13, 16'hff98, 16'hffa4, 16'hff8b, 16'hffc5, 16'hffa6, 16'hffff, 16'h32, 16'hfff7, 16'hffb2, 16'hffb9, 16'hffff, 16'h33, 16'hd, 16'hffd7, 16'hffb0, 16'h23, 16'h88, 16'h24, 16'hffad, 16'hffda, 16'h41, 16'h3a, 16'h5f, 16'h10, 16'hffcf, 16'hffe1, 16'h39, 16'h31, 16'h52, 16'h2e, 16'h17, 16'h11, 16'h73, 16'hffdc, 16'h5, 16'hffc5, 16'hffb9, 16'hffc5, 16'h19, 16'hffcc, 16'hffff, 16'h31, 16'hffcf, 16'hff9f, 16'hffcd, 16'hffea, 16'h25, 16'h33, 16'hffca, 16'hffc3, 16'hffbd, 16'h31, 16'h43, 16'h1b, 16'h3, 16'h36, 16'h1f, 16'h6d, 16'h81, 16'h22, 16'h31, 16'h54, 16'h5e, 16'h4a, 16'h66, 16'h3a, 16'h3c, 16'h38, 16'h46, 16'h1c, 16'h21, 16'hfff1, 16'hd, 16'h32, 16'h67, 16'h28, 16'ha, 16'h6, 16'h8, 16'h16, 16'h15, 16'h22, 16'h2d, 16'h22, 16'hffdc, 16'hfff9, 16'h0, 16'h6, 16'h52, 16'h5a, 16'hc, 16'h23, 16'hfffe, 16'hffff, 16'h46, 16'h2b, 16'h10, 16'h1e, 16'h13, 16'h27, 16'h3e, 16'hf, 16'hffe8, 16'hffea, 16'h11, 16'h1, 16'h21, 16'hffe5, 16'hffcf, 16'hffdd, 16'hffd7, 16'hffb3, 16'hffc0, 16'h2b, 16'h8, 16'hffd3, 16'hffc3, 16'hffbe, 16'hffd6, 16'h33, 16'hffeb, 16'hffcb, 16'hffbb, 16'h20, 16'h2, 16'h17, 16'h1e, 16'h1b, 16'h24, 16'h52, 16'h47, 16'h52, 16'h3e, 16'h3a, 16'h13, 16'h44, 16'h49, 16'h54, 16'h28, 16'h3, 16'h0, 16'hd, 16'hffeb, 16'hffab, 16'hffbe, 16'hffdb, 16'h16, 16'hffde, 16'h8, 16'h56, 16'h73, 16'h3f, 16'h15, 16'hffe1, 16'hffe6, 16'h18, 16'h5d, 16'h88, 16'h49, 16'h5, 16'hff6b, 16'hffd0, 16'h32, 16'h56, 16'h33, 16'hc, 16'hff6b, 16'hff74, 16'hffc7, 16'h28, 16'h20, 16'hfffa, 16'hffc0, 16'hff53, 16'hff7c, 16'hffcf, 16'hffe9, 16'h1c, 16'h5, 16'h3, 16'he, 16'h1f, 16'hf, 16'h26, 16'h14, 16'hffe3, 16'hffcd, 16'hfffc, 16'h25, 16'hff92, 16'hffc7, 16'hffb8, 16'hff8d, 16'hffe5, 16'hffe6, 16'hff1c, 16'hff62, 16'hff71, 16'hff5c, 16'hffa3, 16'hffee, 16'hffb8, 16'hff7a, 16'hff68, 16'hff5e, 16'hffa9, 16'h9, 16'hb, 16'hffda, 16'hffbc, 16'hff9c, 16'hffdc, 16'hfff7, 16'h6, 16'hffe3, 16'hffd4, 16'hff62, 16'hffb4, 16'hb, 16'h10, 16'hffdc, 16'hffe0, 16'hffcc, 16'hffd0, 16'hfff0, 16'h11, 16'h7f, 16'h7f, 16'hfff3, 16'hffc4, 16'hfffe, 16'hffe7, 16'hffee, 16'h1, 16'h31, 16'hffd7, 16'hfff0, 16'hfff3, 16'h48, 16'hd, 16'h40, 16'hfff5, 16'hffaa, 16'h2d, 16'h59, 16'h28, 16'h3c, 16'h15, 16'hffb5, 16'hfff3, 16'h1b, 16'h44, 16'h79, 16'h2f, 16'hffd1, 16'h10, 16'h9, 16'hfffc, 16'hffe6, 16'hff82, 16'hffaa, 16'hfffd, 16'hffea, 16'hff6b, 16'hffe3, 16'hffec, 16'h1b, 16'h12, 16'hfff0, 16'hfeeb, 16'h0, 16'h18, 16'h22, 16'h9, 16'hffe2, 16'hffb2, 16'h33, 16'h23, 16'h5, 16'hffe3, 16'h3, 16'hffd3, 16'h3, 16'h1, 16'h2, 16'h10, 16'hffce, 16'hffbc, 16'hffd6, 16'h5, 16'h1b, 16'hffde, 16'h10, 16'h1f, 16'h2a, 16'hc, 16'h22, 16'h4, 16'h0, 16'h33, 16'h2e, 16'h2, 16'hffdc, 16'h6, 16'h88, 16'h8d, 16'h9e, 16'h38, 16'hffb7, 16'h1, 16'h96, 16'hd9, 16'h10b, 16'h75, 16'hffb4, 16'h12, 16'h92, 16'h10e, 16'h120, 16'h94, 16'hffc5, 16'h32, 16'h2b, 16'h61, 16'h64, 16'h30, 16'hffdb, 16'he, 16'h33, 16'h2d, 16'h7, 16'h15, 16'h17, 16'hffe2, 16'h3, 16'hfffb, 16'ha, 16'h18, 16'hfffc, 16'h12, 16'hffd1, 16'hffbe, 16'hffd3, 16'hffe6, 16'hffd1, 16'h56, 16'h47, 16'h29, 16'hfff5, 16'hffb5, 16'hffa2, 16'h5e, 16'h75, 16'h76, 16'h32, 16'hffe4, 16'hffa7, 16'h14, 16'h4f, 16'h6c, 16'h33, 16'hffe2, 16'hffc9, 16'h1c, 16'hf, 16'hfff2, 16'hffc9, 16'hffa6, 16'hfff3, 16'h1, 16'h34, 16'h48, 16'hffd5, 16'hffb2, 16'hffc3, 16'h1, 16'h70, 16'h64, 16'h30, 16'hffd3, 16'hffde, 16'h21, 16'h76, 16'h6b, 16'h43, 16'hfffa, 16'hffee, 16'hffef, 16'h2d, 16'h3f, 16'h14, 16'hd, 16'hfff8, 16'hffd8, 16'hffe9, 16'h14, 16'hc, 16'h24, 16'h9, 16'hffec, 16'h2c, 16'h36, 16'h1a, 16'h3, 16'ha, 16'hffea, 16'hffef, 16'hc, 16'h4, 16'hffed, 16'hffed, 16'hffe6, 16'hffb9, 16'hffcf, 16'hffed, 16'hffcd, 16'hffd9, 16'hb, 16'h1b, 16'hffe7, 16'h7, 16'hffc9, 16'hffc7, 16'h25, 16'h6b, 16'hc, 16'h29, 16'hffd5, 16'hffd3, 16'hc, 16'h3c, 16'h1d, 16'h12, 16'hffe9, 16'hffdb, 16'hffff, 16'h23, 16'hff89, 16'hff3b, 16'hff99, 16'h7, 16'hfff1, 16'hff96, 16'hffaa, 16'h11, 16'h10, 16'h15, 16'h1, 16'h4e, 16'hffe4, 16'hfff7, 16'ha, 16'h2d, 16'hfff4, 16'h57, 16'h63, 16'h59, 16'h2e, 16'h12, 16'hd, 16'h56, 16'ha1, 16'h82, 16'h52, 16'h25, 16'hfff6, 16'hffb2, 16'hffb7, 16'hffd5, 16'hffd1, 16'hffd0, 16'hffe6, 16'hff7b, 16'h49, 16'h7e, 16'h53, 16'h24, 16'hfff8, 16'hffcf, 16'h1b, 16'h87, 16'hc, 16'hfffe, 16'h65, 16'h2b, 16'hffcf, 16'h71, 16'h1e, 16'h2, 16'h36, 16'h27, 16'hffec, 16'h68, 16'h64, 16'h22, 16'hffc2, 16'hfffb, 16'h12, 16'h43, 16'h69, 16'h2b, 16'hffaf, 16'hffd8, 16'h37, 16'h48, 16'h35, 16'h16, 16'h1, 16'h12, 16'h22, 16'h11, 16'hffd1, 16'hffdd, 16'hffe2, 16'hff75, 16'hff70, 16'hffa8, 16'hffe1, 16'hffc5, 16'h7a, 16'h10a, 16'hbd, 16'h26, 16'h35, 16'h20, 16'h6c, 16'h123, 16'hf5, 16'h38, 16'h1a, 16'h33, 16'h38, 16'h91, 16'h75, 16'hffea, 16'hffd9, 16'hfff3, 16'hffc6, 16'hffb3, 16'hff9e, 16'hff8f, 16'hff9a, 16'hffc9, 16'hfff7, 16'h31, 16'h15, 16'hffaf, 16'hffbc, 16'hffb5, 16'h1a, 16'h30, 16'hffe7, 16'hffac, 16'hffa4, 16'hffdc, 16'hfffb, 16'hab, 16'h84, 16'h7, 16'hffda, 16'h4, 16'hffe1, 16'h2f, 16'h25, 16'h1c, 16'hf, 16'h1a, 16'hfff2, 16'hff9d, 16'hffcb, 16'h25, 16'h7, 16'h24, 16'hfff3, 16'hffd0, 16'hffee, 16'h11, 16'hfff8, 16'hffdf, 16'h9, 16'hffb4, 16'hff4d, 16'hff7c, 16'hffc7, 16'h23, 16'hb, 16'hffd8, 16'hff4b, 16'hff72, 16'hffe4, 16'h40, 16'hffdb, 16'hff61, 16'hff62, 16'hffc4, 16'hffe9, 16'h29, 16'h0, 16'hffaa, 16'hff77, 16'hffc4, 16'hffeb, 16'h54, 16'hfff7, 16'hffbf, 16'hff96, 16'hff99, 16'hffca, 16'h3, 16'hffd1, 16'hff9f, 16'hffa4, 16'hffa0, 16'hffb9, 16'hffd9, 16'hffc5, 16'hff9c, 16'hff74, 16'hff9d, 16'hffcc, 16'h3, 16'h41, 16'h7, 16'hffab, 16'hffd8, 16'hfff4, 16'h26, 16'h8e, 16'ha0, 16'h49, 16'h2b, 16'h1c, 16'h28, 16'h25, 16'h12, 16'hfffd, 16'h12, 16'h37, 16'h3c, 16'hffb5, 16'hffae, 16'hffcd, 16'hfff1, 16'h17, 16'h1e, 16'hfff1, 16'hffa9, 16'hff97, 16'hffc7, 16'hffd4, 16'hffef, 16'h3, 16'h1f, 16'h76, 16'h2a, 16'hf, 16'hffe3, 16'hffdb, 16'hfff5, 16'h3a, 16'h3f, 16'hfff4, 16'hffbc, 16'hfff0, 16'hffee, 16'hffdd, 16'h11, 16'hb, 16'hffea, 16'h6, 16'hffce, 16'hffc3, 16'h2b, 16'h23, 16'h23, 16'h1, 16'hffcf, 16'hfff4, 16'h24, 16'h22, 16'h27, 16'h0, 16'h3f, 16'h3b, 16'h43, 16'h2b, 16'h7, 16'hffeb, 16'hffc8, 16'hff76, 16'hffa4, 16'ha, 16'h3c, 16'h1, 16'hfff9, 16'hffc6, 16'hffdb, 16'h24, 16'h4a, 16'h20, 16'h2c, 16'h50, 16'h42, 16'h47, 16'h3c, 16'hffff, 16'hfffd, 16'h20, 16'h1f, 16'h55, 16'h50, 16'hfff0, 16'hff8b, 16'hffa8, 16'hffd7, 16'hfffd, 16'h5, 16'h7, 16'hffa2, 16'hffd4, 16'hfff3, 16'hffee, 16'hffd6, 16'hfff3, 16'hffdc, 16'hffa2, 16'hffbc, 16'hfff1, 16'h6, 16'hffc7, 16'h3c, 16'ha0, 16'h1f, 16'hffb9, 16'hffcc, 16'hffe0, 16'h40, 16'h5c, 16'hf, 16'hffd2, 16'hffc5, 16'hffcf, 16'hffc9, 16'hffcb, 16'hffb9, 16'hff97, 16'hffc2, 16'hffc4, 16'hff88, 16'hff97, 16'hffb0, 16'hffdf, 16'hffed, 16'hffc2, 16'hffde, 16'hffda, 16'h3, 16'h1a, 16'h7, 16'hfff0, 16'h2d, 16'hffa5, 16'hff7e, 16'hffd3, 16'hffda, 16'h5c, 16'h6d, 16'ha, 16'hff3b, 16'hffaa, 16'hffd2, 16'h6f, 16'h8c, 16'h6f, 16'hff3b, 16'hff62, 16'hffde, 16'hfff0, 16'hfff5, 16'hffbc, 16'hff3d, 16'hff4b, 16'hffbe, 16'hffba, 16'hff88, 16'hff6a, 16'hff37, 16'hff65, 16'hffd3, 16'hffdb, 16'hffc1, 16'hffb6, 16'hff8b, 16'hff86, 16'hffb9, 16'hffe9, 16'hffbb, 16'hffb2, 16'h4, 16'h35, 16'hffe9, 16'hffe6, 16'hff47, 16'hff92, 16'ha1, 16'hb0, 16'h1d, 16'hfffc, 16'h23, 16'h4, 16'h3d, 16'h5a, 16'h2, 16'hffbb, 16'h32, 16'h4e, 16'h34, 16'hfff6, 16'hffd4, 16'hffe9, 16'h31, 16'h1a, 16'h12, 16'hfff0, 16'hffba, 16'hffd7, 16'hb, 16'h46, 16'h53, 16'h32, 16'hfff0, 16'hfffc, 16'hffd1, 16'hffeb, 16'hffda, 16'hc2, 16'ha0, 16'hffbd, 16'hffdb, 16'h27, 16'hffea, 16'h25, 16'h3e, 16'hffef, 16'hffd1, 16'h6, 16'hffb0, 16'h17, 16'h1d, 16'hffce, 16'hff93, 16'hff75, 16'hff9f, 16'hffbc, 16'hffdd, 16'hffd6, 16'hffa5, 16'hffbb, 16'hffc4, 16'hffd3, 16'h6, 16'hfff8, 16'hffb6, 16'hffdf, 16'hffe5, 16'h2, 16'h1b, 16'hffc3, 16'h50, 16'h8e, 16'h31, 16'h14, 16'h1d, 16'hffdd, 16'h18, 16'h4d, 16'h5a, 16'h65, 16'h56, 16'hffcd, 16'ha, 16'h5b, 16'haf, 16'ha7, 16'h4b, 16'hffe5, 16'hc8, 16'hc3, 16'he0, 16'ha1, 16'h1b, 16'hffe4, 16'hc2, 16'hf8, 16'hdd, 16'h6b, 16'h3, 16'hffe0, 16'h23, 16'h63, 16'h58, 16'hf, 16'hffd4, 16'he, 16'h56, 16'h29, 16'h7, 16'h69, 16'h35, 16'hfff9, 16'h30, 16'h3e, 16'h1d, 16'h3a, 16'h10, 16'hffcf, 16'hfff5, 16'h54, 16'h53, 16'h44, 16'h2a, 16'hffca, 16'h10, 16'h58, 16'h5a, 16'h56, 16'h45, 16'hfff0, 16'h32, 16'h25, 16'h27, 16'hfffc, 16'hfff8, 16'hffee, 16'h35, 16'h24, 16'h31, 16'hffee, 16'hffee, 16'h7, 16'hfff3, 16'hffca, 16'h43, 16'h68, 16'h41, 16'hfff6, 16'hff93, 16'hff99, 16'h59, 16'h77, 16'h39, 16'hd, 16'hffc1, 16'hffa0, 16'h68, 16'h7a, 16'h31, 16'h30, 16'h2a, 16'h3, 16'h4, 16'h3, 16'hfff9, 16'h10, 16'h3e, 16'h28, 16'hfffb, 16'hffe9, 16'hffe9, 16'h16, 16'h12, 16'h1, 16'hffef, 16'hffef, 16'h1a, 16'hffe6, 16'h65, 16'h67, 16'hffe8, 16'h38, 16'h51, 16'hffbd, 16'h68, 16'h46, 16'h17, 16'h34, 16'h2d, 16'hffb4, 16'h34, 16'h26, 16'h12, 16'h2, 16'hfff5, 16'hffa4, 16'h10, 16'hffea, 16'hffd4, 16'hffee, 16'h8, 16'hffdd, 16'h8, 16'hffcd, 16'hffc9, 16'hffd7, 16'hfff4, 16'hffc6, 16'h12, 16'hfff0, 16'hfffb, 16'hffe3, 16'hffd4, 16'h25, 16'h1f, 16'hffb5, 16'hff68, 16'hffd6, 16'hfff2, 16'hfffe, 16'hffda, 16'hffbd, 16'hffb4, 16'hffc3, 16'hffd5, 16'hfff1, 16'h42, 16'h52, 16'hf, 16'h1d, 16'hfff6, 16'hffea, 16'h9f, 16'hcf, 16'h84, 16'h1d, 16'he, 16'h4, 16'h91, 16'hc4, 16'ha4, 16'h5d, 16'h19, 16'h0, 16'h55, 16'h7f, 16'h93, 16'h5f, 16'h61, 16'hd, 16'hffc1, 16'h58, 16'hb1, 16'h24, 16'h1c, 16'hffcd, 16'hffaa, 16'h1, 16'h20, 16'hffc5, 16'h19, 16'h49, 16'h17, 16'h44, 16'hff7d, 16'hff6a, 16'h21, 16'hcb, 16'h90, 16'h52, 16'hff87, 16'hff73, 16'hffe6, 16'h70, 16'h46, 16'h9, 16'hff53, 16'hff54, 16'hfff5, 16'h9, 16'hfff3, 16'hff9d, 16'hff4b, 16'hff97, 16'h1, 16'h8, 16'h2d, 16'h15, 16'hf, 16'h19, 16'he, 16'hfff5, 16'hffdb, 16'hff96, 16'hffcd, 16'h16, 16'h41, 16'h4, 16'hff83, 16'hff75, 16'hffa9, 16'hfff9, 16'h18, 16'hffc2, 16'hff9f, 16'hffd6, 16'hb, 16'h1a, 16'hfffa, 16'hffc7, 16'hffb2, 16'hffef, 16'he, 16'h2b, 16'h2a, 16'hfff4, 16'hfff9, 16'h4c, 16'h56, 16'h42, 16'h41, 16'hffe3, 16'h1f, 16'h16, 16'h135, 16'h10d, 16'h40, 16'h5, 16'h24, 16'h22, 16'h99, 16'h76, 16'h12, 16'h28, 16'h9, 16'h43, 16'h14, 16'h17, 16'hffca, 16'h23, 16'hffd1, 16'hffe1, 16'hffb9, 16'hffe0, 16'hffef, 16'h1e, 16'hffb7, 16'hff9a, 16'hffb5, 16'hffc1, 16'hffcf, 16'h1b, 16'hffe1, 16'hffb8, 16'hff8e, 16'hffc7, 16'hffe4, 16'h9, 16'hffac, 16'hff70, 16'hff96, 16'hfff2, 16'hffe4, 16'hfffb, 16'hffd3, 16'hff7c, 16'hffe4, 16'h4b, 16'h22, 16'h22, 16'hffee, 16'hffda, 16'h29, 16'h4a, 16'h16, 16'hfff7, 16'hffb8, 16'hf, 16'h1c, 16'h32, 16'hffee, 16'hf, 16'hffbf, 16'hfff9, 16'hfff0, 16'h19, 16'h21, 16'h12, 16'hffe9, 16'hfff3, 16'hffee, 16'h10, 16'h28, 16'hfffc, 16'hff8c, 16'hffd3, 16'h2e, 16'ha, 16'hfff2, 16'hfff6, 16'hff96, 16'hffae, 16'h11, 16'h7, 16'hfff8, 16'h12, 16'h18, 16'h35, 16'h54, 16'h2b, 16'h13, 16'hffb4, 16'hffe6, 16'h2d, 16'h57, 16'h2b, 16'hc, 16'hffc8, 16'hfffc, 16'he, 16'hffee, 16'hffeb, 16'hfff6, 16'hfff5, 16'hfffd, 16'hffdb, 16'hffd2, 16'hffea, 16'h11, 16'h19, 16'h30, 16'h23, 16'h5f, 16'h3a, 16'h1c, 16'hffeb, 16'h35, 16'h27, 16'h61, 16'h49, 16'h28, 16'hfffb, 16'hffd2, 16'hffe4, 16'h50, 16'h31, 16'h6, 16'hffe7, 16'hff96, 16'hff96, 16'hffff, 16'h0, 16'h0, 16'hffee, 16'hffa9, 16'hffd4, 16'hffe0, 16'hffe5, 16'hfffe, 16'h4, 16'hffec, 16'hffe3, 16'hffe2, 16'hfff2, 16'h1, 16'h10, 16'hffa5, 16'hff75, 16'hfff4, 16'h39, 16'hffe5, 16'h1b, 16'hff8b, 16'hff9c, 16'hffe5, 16'he, 16'hfff1, 16'hffea, 16'h10, 16'h38, 16'hfff2, 16'hfff9, 16'hffe6, 16'hfffc, 16'h2a, 16'h16, 16'hffe5, 16'hfffd, 16'hffd7, 16'hfff6, 16'h23, 16'hffed, 16'hffd4, 16'hffda, 16'hffe9, 16'h10, 16'hfff8, 16'hffc2, 16'hffb4, 16'hffd2, 16'h1, 16'h10, 16'hd, 16'h40, 16'hb, 16'h10, 16'hf, 16'hfff7, 16'hffe5, 16'hffad, 16'hffcd, 16'h2a, 16'h13, 16'h28, 16'hff8e, 16'hff7e, 16'hffde, 16'h44, 16'h13, 16'hffee, 16'hffc2, 16'hffdd, 16'hf, 16'h5f, 16'hfffa, 16'hffef, 16'hffbb, 16'hfff5, 16'hf, 16'h35, 16'hffca, 16'h27, 16'hffad, 16'hff8d, 16'hff7b, 16'hff9a, 16'hffab, 16'hfff1, 16'h28, 16'hff6f, 16'hff8c, 16'hfff9, 16'h30, 16'hffb3, 16'hff89, 16'hff9a, 16'h11, 16'h30, 16'hffef, 16'hff6c, 16'hff48, 16'hffc0, 16'h4e, 16'h17, 16'hfff2, 16'hff97, 16'hffd6, 16'hffdc, 16'h30, 16'hffe7, 16'hffea, 16'hffa6, 16'h27, 16'h4d, 16'haf, 16'h4d, 16'h7, 16'hfff7, 16'h3c, 16'ha6, 16'he0, 16'h56, 16'hfff9, 16'h23, 16'h20, 16'h6d, 16'h1c, 16'hfffb, 16'hd, 16'h0, 16'h110, 16'h142, 16'h9c, 16'h1f, 16'h20, 16'hffe7, 16'h15, 16'h7a, 16'h35, 16'hffee, 16'h25, 16'hffbe, 16'hffa1, 16'hff6f, 16'hff8a, 16'hff88, 16'hffc4, 16'hffd4, 16'hffc1, 16'hff55, 16'hff51, 16'hff7f, 16'hffc1, 16'hffcd, 16'hffbd, 16'hff7a, 16'hff62, 16'hffa1, 16'hffe1, 16'hffeb, 16'h13, 16'h30, 16'hffd0, 16'h97, 16'h60, 16'h1a, 16'hffea, 16'hff89, 16'hfff3, 16'h6d, 16'h75, 16'h9, 16'hc, 16'hff49, 16'hfff4, 16'h5f, 16'h90, 16'hfff9, 16'h3, 16'h28, 16'h45, 16'h17, 16'h7, 16'hfffe, 16'hffdb, 16'h82, 16'h66, 16'h34, 16'h18, 16'h20, 16'h7, 16'h88, 16'h79, 16'h28, 16'hffd0, 16'h22, 16'h61, 16'h8b, 16'h5b, 16'h57, 16'h6e, 16'h6, 16'h48, 16'hb2, 16'h50, 16'h5f, 16'h81, 16'hd, 16'h43, 16'hae, 16'h5b, 16'h12, 16'h2, 16'hffec, 16'hffda, 16'h30, 16'h4, 16'hffd2, 16'hffe5, 16'hfff9, 16'hffba, 16'hff78, 16'hff49, 16'hff8d, 16'hffcd, 16'hfffb, 16'hffd5, 16'hffd6, 16'hffc0, 16'hffbf, 16'hffea, 16'h9, 16'h74, 16'h40, 16'hffce, 16'h48, 16'h31, 16'hffcd, 16'h26, 16'h31, 16'h19, 16'h57, 16'h3f, 16'hffc6, 16'hffa8, 16'hffae, 16'hfff9, 16'h33, 16'h1a, 16'hff98, 16'hffca, 16'hffca, 16'hffda, 16'hffbe, 16'hffe2, 16'hffc7, 16'hffad, 16'hffd7, 16'hffdc, 16'hffb4, 16'hffa7, 16'hffbb, 16'hffdd, 16'hffe6, 16'h3, 16'hfff8, 16'hffc7, 16'hffdc, 16'hffe5, 16'h4a, 16'hfffd, 16'h11, 16'hffd7, 16'hffd0, 16'h49, 16'h6b, 16'hfff6, 16'hfff5, 16'h1, 16'hfff0, 16'h41, 16'h6b, 16'h39, 16'h10, 16'h24, 16'hfffd, 16'h32, 16'h1b, 16'h15, 16'hffea, 16'h19, 16'hfffc, 16'hb, 16'h20, 16'h9, 16'h6, 16'h3e, 16'hffd3, 16'hffe8, 16'h17, 16'ha, 16'ha, 16'h4, 16'h15, 16'h71, 16'h7e, 16'hfff0, 16'h35, 16'h3c, 16'h21, 16'h16, 16'h25, 16'h35, 16'h67, 16'h65, 16'hffeb, 16'hff85, 16'hff88, 16'hffc3, 16'hffd7, 16'hffe9, 16'hffe8, 16'hff9c, 16'hffc4, 16'hffd7, 16'hffd2, 16'hffb7, 16'hffee, 16'hffac, 16'hfff8, 16'hffe8, 16'hfff5, 16'hffc2, 16'h1, 16'hfff6, 16'h37, 16'h38, 16'h2d, 16'hffef, 16'hffed, 16'hffe0, 16'h122, 16'h121, 16'h73, 16'hffcc, 16'hffc4, 16'hd5, 16'h100, 16'h91, 16'h7f, 16'hffeb, 16'hffc8, 16'h94, 16'hc7, 16'ha2, 16'h87, 16'h15, 16'hfff5, 16'h8f, 16'hd0, 16'hb6, 16'h87, 16'h14, 16'hffe2, 16'h7e, 16'hbe, 16'h99, 16'h56, 16'h24, 16'hffc0, 16'h60, 16'h81, 16'h7a, 16'h34, 16'h11, 16'h2f, 16'ha5, 16'hfffe, 16'hffa3, 16'hffb2, 16'hffc1, 16'h7f, 16'h8b, 16'h12, 16'hff74, 16'hffb2, 16'hffc4, 16'h21, 16'h24, 16'h13, 16'hff72, 16'hff9e, 16'hffcf, 16'h2f, 16'h1a, 16'hfff2, 16'hff8b, 16'hff8a, 16'hffc9, 16'h44, 16'h2d, 16'h20, 16'hffa3, 16'hffc1, 16'hffbd, 16'h65, 16'h35, 16'h36, 16'hfff3, 16'hffdd, 16'hffd7, 16'hfffa, 16'hffba, 16'hff9f, 16'hffcc, 16'hffb5, 16'hffd7, 16'h2b, 16'hffed, 16'hffc9, 16'hffa8, 16'hffc8, 16'hffea, 16'hfffa, 16'hff79, 16'hff48, 16'hff6c, 16'hff93, 16'hffdd, 16'hffcd, 16'hff48, 16'hff62, 16'hffab, 16'hffde, 16'hfff4, 16'h15, 16'hffe9, 16'hffe1, 16'h0, 16'h12, 16'hffe9, 16'hfff9, 16'hfffc, 16'h2b, 16'h35, 16'h16, 16'h8, 16'hffbe, 16'hffd2, 16'hffd1, 16'h26, 16'h1d, 16'h1e, 16'hffe3, 16'hffbb, 16'hffae, 16'hfff6, 16'hb, 16'h2c, 16'hffc1, 16'hff99, 16'hff8f, 16'hffcd, 16'hffed, 16'hc, 16'hfff4, 16'hffd1, 16'hffd8, 16'hffd7, 16'h1, 16'h22, 16'hffd1, 16'hffe2, 16'hffcc, 16'hffc1, 16'hffe0, 16'h23, 16'hfff2, 16'hffd8, 16'hfff0, 16'hffeb, 16'h16, 16'h57, 16'hffb9, 16'h4b, 16'h49, 16'h22, 16'hffeb, 16'hfff3, 16'hffdb, 16'h6, 16'h1b, 16'hffef, 16'hffcc, 16'hffe1, 16'hffde, 16'hfffe, 16'hffdf, 16'hffec, 16'hffc9, 16'hfff8, 16'hffda, 16'hffb4, 16'hff99, 16'hffc2, 16'hffe0, 16'hfff8, 16'hffd5, 16'hffed, 16'hffe2, 16'hffe3, 16'h10, 16'h6, 16'hffea, 16'hfffc, 16'h50, 16'h4a, 16'h5f, 16'hffe4, 16'h53, 16'h8c, 16'h95, 16'h5b, 16'h35, 16'h19, 16'hfffd, 16'h3a, 16'h30, 16'h12, 16'h22, 16'hfffc, 16'h18, 16'hffee, 16'hffe4, 16'hffcf, 16'hfffc, 16'hffff, 16'h19, 16'hffe9, 16'hffea, 16'hfffb, 16'h4, 16'h18, 16'h2e, 16'h21, 16'h1b, 16'h31, 16'h36, 16'h2f, 16'h17, 16'h4e, 16'h41, 16'h5b, 16'h69, 16'h44, 16'h22, 16'hffc1, 16'hff53, 16'hff8f, 16'hffa3, 16'h13, 16'h4f, 16'hffb0, 16'hff6e, 16'hff9b, 16'hffb9, 16'hfff3, 16'h3d, 16'hffea, 16'hffc4, 16'hff8c, 16'hffb0, 16'hfff9, 16'h38, 16'hffcd, 16'hffd5, 16'hffca, 16'hffd4, 16'hffdb, 16'h10, 16'hffb8, 16'hffd0, 16'hffc5, 16'hffd9, 16'hffec, 16'h16, 16'hffe1, 16'hffbb, 16'hffbd, 16'hffe1, 16'hfff3, 16'hffce, 16'h86, 16'h79, 16'h15, 16'hfff7, 16'h36, 16'hffcb, 16'h49, 16'h13, 16'hffcc, 16'hffcb, 16'h1e, 16'hffcb, 16'hfffd, 16'ha, 16'hfff9, 16'hfff0, 16'h1c, 16'hffee, 16'h14, 16'hfff3, 16'h3, 16'h10, 16'h1e, 16'hfffd, 16'h29, 16'h4, 16'h2b, 16'h26, 16'h23, 16'hfff3, 16'h4f, 16'h35, 16'h62, 16'h56, 16'h45, 16'h1e, 16'h21, 16'h37, 16'h93, 16'h68, 16'h2a, 16'h1e, 16'h34, 16'ha5, 16'h71, 16'h46, 16'hffee, 16'he, 16'h78, 16'h79, 16'h4d, 16'h2c, 16'hfffb, 16'h29, 16'h4b, 16'h1c, 16'hb, 16'h17, 16'hfff7, 16'h25, 16'hffc2, 16'hffd3, 16'hffc6, 16'hffb5, 16'hfffd, 16'h1d, 16'h3, 16'hffa0, 16'hff63, 16'hff79, 16'he, 16'h6, 16'h1b, 16'h17, 16'hffe9, 16'hffe3, 16'h30, 16'h3f, 16'h60, 16'h18, 16'hffbd, 16'h15, 16'h2b, 16'h78, 16'h6f, 16'h11, 16'h23, 16'h22, 16'h1, 16'hfff5, 16'hffc1, 16'hfff1, 16'h4a, 16'h6d, 16'h19, 16'hffb0, 16'hffc0, 16'h57, 16'hc1, 16'hf4, 16'h42, 16'hffda, 16'hfffc, 16'hb7, 16'h119, 16'h11a, 16'h42, 16'h15, 16'hd, 16'h2, 16'h13, 16'hfff5, 16'h3a, 16'h1b, 16'hff9a, 16'hff67, 16'hffb3, 16'hffe7, 16'h25, 16'h20, 16'h41, 16'h67, 16'h6e, 16'hfffa, 16'hffe6, 16'hffdd, 16'hffeb, 16'h26, 16'h60, 16'h15, 16'h6, 16'hc, 16'hffb3, 16'hffbc, 16'hffb4, 16'hffc4, 16'h1b, 16'h27, 16'hffbc, 16'hff78, 16'hff4e, 16'hff85, 16'ha, 16'h1f, 16'h44, 16'hf, 16'h3, 16'hffeb, 16'hfff2, 16'hfffb, 16'h30, 16'hffec, 16'h24, 16'hfffa, 16'hffe8, 16'h3a, 16'hffc4, 16'hffbf, 16'h22, 16'hfffc, 16'hffaa, 16'h3e, 16'hff95, 16'hff58, 16'hffde, 16'hffe2, 16'hffcf, 16'h2e, 16'hffd5, 16'hff8a, 16'h2d, 16'h1b, 16'h23, 16'hc, 16'h8, 16'h29, 16'h8f, 16'h62, 16'h43, 16'h14, 16'h8, 16'h2e, 16'h57, 16'h14, 16'hb, 16'h12, 16'h37, 16'h2d, 16'h20, 16'hffe9, 16'hffb0, 16'h11, 16'hffb2, 16'hff82, 16'hffe3, 16'hffd1, 16'hff99, 16'hfff3, 16'hffbb, 16'hff99, 16'hffab, 16'hffac, 16'hffb5, 16'ha, 16'hffa8, 16'hff99, 16'hff6b, 16'hff9a, 16'h8, 16'hfff5, 16'hffd0, 16'hffe8, 16'hffd4, 16'hffed, 16'h23, 16'h0, 16'hffe5, 16'h26, 16'h48, 16'h13, 16'hffe5, 16'h2f, 16'h36, 16'h2f, 16'hc, 16'h3, 16'hffb5, 16'hffd7, 16'h21, 16'hffdf, 16'hffc0, 16'hffaa, 16'hff96, 16'hffc4, 16'hffb4, 16'hffa0, 16'hffe9, 16'hffe3, 16'hffc3, 16'hffe2, 16'hff6d, 16'hff86, 16'hffdc, 16'h1d, 16'h1, 16'hffea, 16'hffb2, 16'hffce, 16'hfff3, 16'h36, 16'h44, 16'hffdf, 16'h1, 16'hffc8, 16'hffc2, 16'hffaa, 16'hffdd, 16'hc, 16'hffd4, 16'hff8c, 16'hff5d, 16'hffb4, 16'hffff, 16'hffe8, 16'hffb1, 16'hffb7, 16'hffc4, 16'hffcb, 16'hffef, 16'hfff1, 16'hfff9, 16'hffe4, 16'hffef, 16'hffde, 16'hffe7, 16'hfff3, 16'h5b, 16'h31, 16'he, 16'hffeb, 16'hfff8, 16'h1e, 16'h13, 16'h29, 16'h20, 16'h17, 16'hfff0, 16'h34, 16'hffc4, 16'h11, 16'h3e, 16'hf, 16'hb, 16'h29, 16'h2a, 16'h28, 16'h10, 16'hffde, 16'hffd4, 16'h5, 16'h28, 16'h2a, 16'hfffd, 16'hfff1, 16'hffe5, 16'hfffd, 16'hffcb, 16'hffc8, 16'hffe8, 16'h2f, 16'h13, 16'hfffb, 16'hff9e, 16'hffc7, 16'h17, 16'h4b, 16'h37, 16'hf, 16'hffc5, 16'h3b, 16'h85, 16'h74, 16'h67};
    // logic signed [15:0] threshold [0:OC-1] = {-16'd31, -16'd73, -16'd16, -16'd33, -16'd13, -16'd3, -16'd1543, -16'd4, -16'd8, -16'd14};
    logic [CONV1_IMG_OUT_SIZE*CONV1_IMG_OUT_SIZE-1:0] conv1_img_out [0:CONV1_OC-1];
    logic [POOL1_IMG_OUT_SIZE*POOL1_IMG_OUT_SIZE-1:0] pool1_img_out [0:CONV1_OC-1];
    logic [CONV2_IMG_OUT_SIZE*CONV2_IMG_OUT_SIZE-1:0] conv2_img_out [0:CONV2_OC-1];
    logic [POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE-1:0] pool2_img_out [0:CONV2_OC-1];
    logic [FC_IC-1:0] fc_in;
    logic signed [15:0] fc_out [0:FC_OC-1];
    logic [OUTPUT_BIT-1:0] result;

    Conv2d #(
        .IC(CONV1_IC),
        .OC(CONV1_OC),
        .IMG_IN_SIZE(CONV1_IMG_IN_SIZE)
    ) conv1 (
        .img_in(conv1_img_in),
        .weights(conv1_weights),
        // .threshold(threshold),
        .img_out(conv1_img_out)
    );

    MaxPool2d #(
        .IC(CONV1_OC),
        .IMG_IN_SIZE(CONV1_IMG_OUT_SIZE)
    ) pool1 (
        .img_in(conv1_img_out),
        .img_out(pool1_img_out)
    );

    Conv2d #(
        .IC(CONV1_OC),
        .OC(CONV2_OC),
        .IMG_IN_SIZE(POOL1_IMG_OUT_SIZE)
    ) conv2 (
        .img_in(pool1_img_out),
        .weights(conv2_weights),
        // .threshold(threshold),
        .img_out(conv2_img_out)
    );

    MaxPool2d #(
        .IC(CONV2_OC),
        .IMG_IN_SIZE(CONV2_IMG_OUT_SIZE)
    ) pool2 (
        .img_in(conv2_img_out),
        .img_out(pool2_img_out)
    );

    genvar conv2_oc;
    generate
        for (conv2_oc=0; conv2_oc<CONV2_OC; conv2_oc=conv2_oc+1) begin
            assign fc_in[conv2_oc*POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE +: POOL2_IMG_OUT_SIZE*POOL2_IMG_OUT_SIZE] = pool2_img_out[conv2_oc];
        end
    endgenerate

    FC #(
        .IC(FC_IC),
        .OC(FC_OC)
    ) fc (
        .in(fc_in),
        .weights(fc_weights),
        .out(fc_out)
    );

    Comparator #(
        .IC(FC_OC),
    ) compare (
        .in(fc_out),
        .out(result)
    );

    wire _unused_ok = &{result};

endmodule

