`timescale 1ns/1ps
`include "bnn_network.sv"

module toplayer();

    parameter int IMG_SIZE = 30;
    parameter int BNN1_CHANL = 8;
    parameter int BNN2_CHANL = 16;
    parameter int KERNEL_SIZE = 3;
    parameter int MAXPOOL_KERNEL_SIZE = 2;
    parameter int MAXPOOL_STRIDE = 2;
    parameter int MLP_CHANL = 32;
    parameter int NUM_CLASS = 10;
    parameter int DEFAULT_THRESHOLD_WIDTH = 8;

    parameter int BNN1_IMG_SIZE = IMG_SIZE-KERNEL_SIZE+1;
    parameter int MAXPOOL1_IMG_SIZE = BNN1_IMG_SIZE/MAXPOOL_STRIDE;
    parameter int BNN2_IMG_SIZE = MAXPOOL1_IMG_SIZE-KERNEL_SIZE+1;
    parameter int MAXPOOL2_IMG_SIZE = BNN2_IMG_SIZE/MAXPOOL_STRIDE;

    logic [IMG_SIZE*IMG_SIZE-1:0] img;
    logic [KERNEL_SIZE*KERNEL_SIZE*BNN1_CHANL] bnn1_weights;
    logic [KERNEL_SIZE*KERNEL_SIZE*BNN1_CHANL*BNN2_CHANL] bnn2_weights;
    logic [BNN2_CHANL*MAXPOOL2_IMG_SIZE*MAXPOOL2_IMG_SIZE*MLP_CHANL] mlp1_weights;
    logic [MLP_CHANL*NUM_CLASS] mlp2_weights;
    logic [31:0] bnn1_threshold;
    logic [111:0] bnn2_threshold;
    logic [319:0] mlp1_threshold;
    logic [$clog2(NUM_CLASS)-1:0] out;
    
    
    assign img = 'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000011111110000000000000000000000111111111000000000000000000001111000111000000000000000000011110000011100000000000000000011100000011100000000000000000011100000011100000000000000000011100000011100000000000000000011100000011100000000000000000011100000011100000000000000000001100000011100000000000000000001110000011000000000000000000001110000111000000000000000000001110001110000000000000000000000111111110000000000000000000000111111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign bnn1_weights = 'h1900B80377DC07F3F6;
    assign bnn2_weights = 'h8DFEE00FF07FFE070F4EC025A647F803FCF72BD53EE3FD9F2765BFDFB7D7EC17901865BE58C974C06DB88BA7D71100081FFCAD1BFC417338AE2EDFE89A7FBBAE0926CF3DFEFF7729110FFFD03E12F3C1D8B48092700F5A07FFFAF871E3FC03C75C703BBA43D5326E3C02FDF7FCB1869B32FA00FB7F3BEDBEE076FA6996F7C6EBA9C606DC99B2EB3CDBAB6E7DB763A5B7;
    assign mlp1_weights = 'h3FFBFFFFFE7C8825C364EFBAE14F5F7ADBD405BFF410318584300FA452FB8608011DDDBE2FAC7FFCFCD251307A7BEFFFFDD97CBC7B960FDC033AF6DDFFFC18EDA638A9B69EDFFF4EC208308166FE946BEA359511FD85CF3CFBA1BC4E300B43C73E384F7FF3DEFD1AF8031609B3BE9EF8EF3E1038AAE3E53C33E32D138DC71011F81FF2C2228E3DB38629BCF03A9905E1149E51C5968F10117BC64C74798EBEC6189F7240407FA1831CEF9C226B86FCCD475AD708EBFED122E86E0006B0EBA6DC0C3B5942073DE400E0B687B020E7FFDFF1001B8FC9138EB764FF9E764166411C6328FF7DE16980270C72ABCE3B643E77F93A8171F619C0101A738C009AAA3057AB5A6E1C83909E69779947EB3663ADDCB1C835EC719EC341D2B9E5F836FBE671B30820C096775CFFBE2A6085FFF847BBFD952D7DC7BFC0287208399B75CFBBCE5C140CF81D290A13CBBCF2C7BB0E39023BA3D485F7B810108DF38E66BC13BC56F04FDF89D59473BE8C46002505E573E7FCF0E03A9C79DD9AD59F766BD1BF2C04ADA53036B7F72F4DDBADD37F19F7E6F307BECD8EECDFB58942182613E13C7A28CCF70C8F9A493C106130CE0D1A0A6557BE70C1821CD800037A1201004EEEEBEF7F1BE078000AA04AA384E9818B9E7B138FAE8B45ADFADFE9DBA8248ADF7CF3DE001530000F500D18107F4227100812E66000EA66C51A02D67CF3B11E74015E0009AB38B83B3E5D1A1B2B4448100080679CF7F84418020001DFC5EFCEAF1C837FF0B2974C23461018A60ECB4C0D1AD9F1891AE851ED0410BAE63C60AC61FD283AC2890872F8E75FF2E9EF44EFEC4D3F27FF2B015E7C6B6343863C433A71E185F26052AFA0138800E09EF5FFBA8DE2863CACEBA75FF458ECBBDF3F0C498302281CBBB61F21E66DC62EC83060010D5800CBDFEC80605133E03BE7B5FFF4214507F779F25FC9EFBF7D01EFFE4B5E5FFFDF782DF80605CF7DF3FEB34EBC5197C71E5B1DB7F237BA4679C422108C478458045CF9FDCFF50308041D37714104F7AD106164E5D9101673FE80000AE2C300AF7BFBCE15FE001DFFFF5A9C18038AA4BFF7FFFBFF68404459B0206C4206D714FFC4C388028459831E7FA4FCFFFF6EB5B024F104FA465FFE9C91222E9E9B1ECF2E1438600518810801B6F590ED98214C1CF081EF20C3A8301E39FFF97970B3B9F59C0F87C007AA7FF5ED9F1AC80C3A0095BCF28071E384447DF5D7C34FB100048A0EA401867FF2C24CFCB9F1EF0FEDCFFD75C4F76C34FE2FF7CF5C41EE705792FEF0C08003AD00C7CF8FBE1418F5FF9C11D2C1B41A407EB31010C5C7133F74AEF0FEFBCCA53AFA6D4F2C651C8BEFBEFF0CDF39FD4A1EFAFE74B0FC31A5F7396388734265F2DDF96D800871C7367AEB7585C3FBF68697FFFFF3DD5759C1F3DEF9CDF977F277DFFBFE0D0915BDA4903EEFBE1C7F9851ED91C5436002003020F6102420065106FF5B67FFFB70841B09F12D7FFFFFFFFE3F2A69C3E1811533DF9B2C3F17698204A1F77FD3FF1FEBFFFF3F318063FBC18B2BDAFF94E2078AAF1ECF7FFC30026109D078C030AE738AE3CDC034F1B04379F4E1F7D315F9A7D7B966D7FFFE0A2CDD18308BF7CFF738587FBC51A4F5C3F28E0C61860EB81F28F3E8E86B6FD77D2C75E6FFB0756B36734DFFDF6197BF7B760B19B4C6FD9809ED6F384F4940EE0861D327192927F7F6209249FE165A75F3D520808B07BE9106E75B7C800E0506C3FFF91073013C25A20C4200B75D98F28F3CFFFFF97C1C156067A5FCC127B6003001F325CBDB15800004000D219FDFCC3E418C276A83EB82408278AE3477A511536BF38C3EF1C9041E29057305FEFF990CF8144C820235F0FB241800A1A6E1E283AA08234FD2E10628023C140968AD478E309369456FBC5811005AF00EF38F0D0F7547E71FDE09A5AE27C6080038F4DF33C75663F007BCAAB96FE394E3C84063FF4FDDFD5E7DFB8002281ADC77DF21EB003C0D46548F4FE59000000F6F87576E98E79F78F0C9A0021445B8D9AE638DD483CC0A2804A47DEC6DF6B8DE610D31370C79C2705BFB0861CEC9A320B058E3CD6396C715D6D8A2D28CE73F30F997B0D8620C30D366358F3891D219C20CE618C630FE12B2029FAE98C7BB7BFFE100790182B0407B8F7607EAA30009769E08BDA410F2DDEF90861C3B28C7DED69420C90C413DAB80D10C1097BDF30620A025D0E820561290A373FBF706259A7C1491C2EA000006C7A7654F7F1EBD5B4FB3AE88CBBFC0008F6592EBDECF80A7EF5CFDFC1062FC64E7F56ADBE681862E1FED753163CE018F1E3A4C327323987F1CBFFA5C7DE7E3C51FF78EFD4778B3E7C018FC914E1DFF6825C45DFF83A7FF247F5CC95B7BE9B10078713B7861D6D7180B7BEB104601038FBF8BFBD9328C025F71267E7F3D20F1DFE20BF8049F9EBCFAC746FBF720EFFC8A9C70C7A8BC06014737ACFEBA6339BA4AD0611E088913C79EE7AF78FBFE629649C37F3A458C32DDC4CE180813438E3FF59E394E04C36C99003EFD982F2FDB89F43E6A9A382BBCE7FBEFF1063F5D1F643F53C99DFF87F2AA1C98F079FFFA55931FEFDF891479FFF5B9FDD681EF752386C56C1AC848F386C104721D9C6E307CFEDD06161FBFD1DDDEFE00897F1BDD7B47BBFFBE7C89230BE5583722BF3954AB12182E0C6E39228824C41022C0180055B7D505FB87EA19D4855B429AD000529F410E30899BEA04226110E51491BB0E3339258AA440B31ABE8ABBF348007102F880029264C80814828437FB187E18880982EFDFCEA43050C513BEE830CA9E61A17BF8B4F83AF0801000001003229F05367FE63CE002E70000CBFD92D10542C08008BEB0F9DDDE7AF804A2EBE2910B773DDFE3D7EFFFC101E6DDE9C11E65B77D042CE79F11CEE731FE3E401D7085961EFFF145B67FF0519EDD2E67FDFEBFDC7093AD860803AEDF2D08AF8877E30C2FA06FFAE5FE0BB7BF20D88018155473FFFF2238E19F78F300277DEB64B5F5E0BC78021CD3F423FFF99C38638D4F5C6BBD61D547EFC702467DFFE74FF6417FD78118FFE2F9F3BFBA58533FF0260BFAFEF0B79AE352957577FF78A101021A1282086093EDE2FE71C1E1ECF762E1317DE6907DF7FF4764BB0F6F282ADDFD800603FFF29E78BCB0FFE70DFDFF87500022200E40FAFE5F883CFB5C9DD038F7C4D87FFF7E14D6A600F62121AF7FFB7DF3F821B201CFA21BF67FEA62A468BA7A90E39BEC182707AD021C17E3FFE43F6A67C708E4B7DF51;
    assign mlp2_weights = 'h0C9D7B772330FCB0B03727E6ECE239C3B115C4FF8E7F082F2E794C77A76A96FA6E4CDACD50495098;
    assign bnn1_threshold = 'h45454546;
    assign bnn2_threshold = 'h0810204081420408183040810205;
    assign mlp1_threshold = 'h48120481204812048120481204812048120481204812048120481204812048120481204812048120;
    
    BNN_network netowrk (
        .in_image(img),
        .bnn1_weights(bnn1_weights),
        .bnn2_weights(bnn2_weights),
        .mlp1_weights(mlp1_weights),
        .mlp2_weights(mlp2_weights),
        .bnn1_threshold(bnn1_threshold),
        .bnn2_threshold(bnn2_threshold),
        .mlp1_threshold(mlp1_threshold),
        .out(out)
    );

endmodule


module tb_toplayer();

  // Instantiate your DUT (toplayer)
  toplayer dut();

  // Generate a dummy clock signal to force time progression.
  logic clk;
  initial begin
    clk = 0;
    forever #5 clk = ~clk;  // 10 ns period clock.
  end

  // Dummy sequential process to ensure clock is used.
  logic dummy_reg;
  always_ff @(posedge clk) begin
    dummy_reg <= ~dummy_reg;
  end

  // Dump waveforms for viewing
  initial begin
    $dumpfile("tb_toplayer.vcd");
    $dumpvars(0, tb_toplayer);
  end

  // Stimulus: Wait a while, print outputs, then finish simulation.
  initial begin
    // Wait for a few clock cycles (say 100 ns).
    #100;
    $display("Simulation Time: %0t ns", $time);
    $display("Image: %b", dut.img);
    $display("BNN Network Output: %h", dut.out);
    #10;
    $finish;
  end

endmodule