module MLP_Neuron #(

)(
    input wire []
);


endmodule